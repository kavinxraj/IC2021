/*********************************************************/
// MODULE: 
//
// FILE NAME: dum.sv 
// VERSION: 0.1
// DATE: 2021-Sep-20 
// AUTHOR: KavinRaj D
//
// CODE TYPE: RTL or Behavioral Level
//
// DESCRIPTION:
//
/*********************************************************/

module dum
(
	input x,
	output logic y
);

assign y = x;

endmodule
