module csa
#(
	parameter DEPTH = 63,
	parameter WIDTH = 6
)
(
	input [DEPTH-1:0] i,
	output [WIDTH-2:0] sum,
	output cy
);
localparam MAX_STAGES = WIDTH;

logic [MAX_STAGES-1:0][DEPTH:0] s,c;		//Number of Wires not accurate

csa3 csa_s0_a0(
					.a( i[0] ),
					.b( i[1] ),
					.c( i[2] ),
					.sum( s[0][0] ),
					.cy( c[0][0] ));
csa3 csa_s0_a1(
					.a( s[0][0] ),
					.b( i[3] ),
					.c( i[4] ),
					.sum( s[0][1] ),
					.cy( c[0][1] ));
csa3 csa_s0_a2(
					.a( s[0][1] ),
					.b( i[5] ),
					.c( i[6] ),
					.sum( s[0][2] ),
					.cy( c[0][2] ));
csa3 csa_s0_a3(
					.a( s[0][2] ),
					.b( i[7] ),
					.c( i[8] ),
					.sum( s[0][3] ),
					.cy( c[0][3] ));
csa3 csa_s0_a4(
					.a( s[0][3] ),
					.b( i[9] ),
					.c( i[10] ),
					.sum( s[0][4] ),
					.cy( c[0][4] ));
csa3 csa_s0_a5(
					.a( s[0][4] ),
					.b( i[11] ),
					.c( i[12] ),
					.sum( s[0][5] ),
					.cy( c[0][5] ));
csa3 csa_s0_a6(
					.a( s[0][5] ),
					.b( i[13] ),
					.c( i[14] ),
					.sum( s[0][6] ),
					.cy( c[0][6] ));
csa3 csa_s0_a7(
					.a( s[0][6] ),
					.b( i[15] ),
					.c( i[16] ),
					.sum( s[0][7] ),
					.cy( c[0][7] ));
csa3 csa_s0_a8(
					.a( s[0][7] ),
					.b( i[17] ),
					.c( i[18] ),
					.sum( s[0][8] ),
					.cy( c[0][8] ));
csa3 csa_s0_a9(
					.a( s[0][8] ),
					.b( i[19] ),
					.c( i[20] ),
					.sum( s[0][9] ),
					.cy( c[0][9] ));
csa3 csa_s0_a10(
					.a( s[0][9] ),
					.b( i[21] ),
					.c( i[22] ),
					.sum( s[0][10] ),
					.cy( c[0][10] ));
csa3 csa_s0_a11(
					.a( s[0][10] ),
					.b( i[23] ),
					.c( i[24] ),
					.sum( s[0][11] ),
					.cy( c[0][11] ));
csa3 csa_s0_a12(
					.a( s[0][11] ),
					.b( i[25] ),
					.c( i[26] ),
					.sum( s[0][12] ),
					.cy( c[0][12] ));
csa3 csa_s0_a13(
					.a( s[0][12] ),
					.b( i[27] ),
					.c( i[28] ),
					.sum( s[0][13] ),
					.cy( c[0][13] ));
csa3 csa_s0_a14(
					.a( s[0][13] ),
					.b( i[29] ),
					.c( i[30] ),
					.sum( s[0][14] ),
					.cy( c[0][14] ));
csa3 csa_s0_a15(
					.a( s[0][14] ),
					.b( i[31] ),
					.c( i[32] ),
					.sum( s[0][15] ),
					.cy( c[0][15] ));
csa3 csa_s0_a16(
					.a( s[0][15] ),
					.b( i[33] ),
					.c( i[34] ),
					.sum( s[0][16] ),
					.cy( c[0][16] ));
csa3 csa_s0_a17(
					.a( s[0][16] ),
					.b( i[35] ),
					.c( i[36] ),
					.sum( s[0][17] ),
					.cy( c[0][17] ));
csa3 csa_s0_a18(
					.a( s[0][17] ),
					.b( i[37] ),
					.c( i[38] ),
					.sum( s[0][18] ),
					.cy( c[0][18] ));
csa3 csa_s0_a19(
					.a( s[0][18] ),
					.b( i[39] ),
					.c( i[40] ),
					.sum( s[0][19] ),
					.cy( c[0][19] ));
csa3 csa_s0_a20(
					.a( s[0][19] ),
					.b( i[41] ),
					.c( i[42] ),
					.sum( s[0][20] ),
					.cy( c[0][20] ));
csa3 csa_s0_a21(
					.a( s[0][20] ),
					.b( i[43] ),
					.c( i[44] ),
					.sum( s[0][21] ),
					.cy( c[0][21] ));
csa3 csa_s0_a22(
					.a( s[0][21] ),
					.b( i[45] ),
					.c( i[46] ),
					.sum( s[0][22] ),
					.cy( c[0][22] ));
csa3 csa_s0_a23(
					.a( s[0][22] ),
					.b( i[47] ),
					.c( i[48] ),
					.sum( s[0][23] ),
					.cy( c[0][23] ));
csa3 csa_s0_a24(
					.a( s[0][23] ),
					.b( i[49] ),
					.c( i[50] ),
					.sum( s[0][24] ),
					.cy( c[0][24] ));
csa3 csa_s0_a25(
					.a( s[0][24] ),
					.b( i[51] ),
					.c( i[52] ),
					.sum( s[0][25] ),
					.cy( c[0][25] ));
csa3 csa_s0_a26(
					.a( s[0][25] ),
					.b( i[53] ),
					.c( i[54] ),
					.sum( s[0][26] ),
					.cy( c[0][26] ));
csa3 csa_s0_a27(
					.a( s[0][26] ),
					.b( i[55] ),
					.c( i[56] ),
					.sum( s[0][27] ),
					.cy( c[0][27] ));
csa3 csa_s0_a28(
					.a( s[0][27] ),
					.b( i[57] ),
					.c( i[58] ),
					.sum( s[0][28] ),
					.cy( c[0][28] ));
csa3 csa_s0_a29(
					.a( s[0][28] ),
					.b( i[59] ),
					.c( i[60] ),
					.sum( s[0][29] ),
					.cy( c[0][29] ));
csa3 csa_s0_a30(
					.a( s[0][29] ),
					.b( i[61] ),
					.c( i[62] ),
					.sum( s[0][30] ),
					.cy( c[0][30] ));
assign sum[0] = s[0][30];

csa3 csa_s1_a0(
					.a( c[0][0] ),
					.b( c[0][1] ),
					.c( c[0][2] ),
					.sum( s[1][0] ),
					.cy( c[1][0] ));
csa3 csa_s1_a1(
					.a( s[1][0] ),
					.b( c[0][3] ),
					.c( c[0][4] ),
					.sum( s[1][1] ),
					.cy( c[1][1] ));
csa3 csa_s1_a2(
					.a( s[1][1] ),
					.b( c[0][5] ),
					.c( c[0][6] ),
					.sum( s[1][2] ),
					.cy( c[1][2] ));
csa3 csa_s1_a3(
					.a( s[1][2] ),
					.b( c[0][7] ),
					.c( c[0][8] ),
					.sum( s[1][3] ),
					.cy( c[1][3] ));
csa3 csa_s1_a4(
					.a( s[1][3] ),
					.b( c[0][9] ),
					.c( c[0][10] ),
					.sum( s[1][4] ),
					.cy( c[1][4] ));
csa3 csa_s1_a5(
					.a( s[1][4] ),
					.b( c[0][11] ),
					.c( c[0][12] ),
					.sum( s[1][5] ),
					.cy( c[1][5] ));
csa3 csa_s1_a6(
					.a( s[1][5] ),
					.b( c[0][13] ),
					.c( c[0][14] ),
					.sum( s[1][6] ),
					.cy( c[1][6] ));
csa3 csa_s1_a7(
					.a( s[1][6] ),
					.b( c[0][15] ),
					.c( c[0][16] ),
					.sum( s[1][7] ),
					.cy( c[1][7] ));
csa3 csa_s1_a8(
					.a( s[1][7] ),
					.b( c[0][17] ),
					.c( c[0][18] ),
					.sum( s[1][8] ),
					.cy( c[1][8] ));
csa3 csa_s1_a9(
					.a( s[1][8] ),
					.b( c[0][19] ),
					.c( c[0][20] ),
					.sum( s[1][9] ),
					.cy( c[1][9] ));
csa3 csa_s1_a10(
					.a( s[1][9] ),
					.b( c[0][21] ),
					.c( c[0][22] ),
					.sum( s[1][10] ),
					.cy( c[1][10] ));
csa3 csa_s1_a11(
					.a( s[1][10] ),
					.b( c[0][23] ),
					.c( c[0][24] ),
					.sum( s[1][11] ),
					.cy( c[1][11] ));
csa3 csa_s1_a12(
					.a( s[1][11] ),
					.b( c[0][25] ),
					.c( c[0][26] ),
					.sum( s[1][12] ),
					.cy( c[1][12] ));
csa3 csa_s1_a13(
					.a( s[1][12] ),
					.b( c[0][27] ),
					.c( c[0][28] ),
					.sum( s[1][13] ),
					.cy( c[1][13] ));
csa3 csa_s1_a14(
					.a( s[1][13] ),
					.b( c[0][29] ),
					.c( c[0][30] ),
					.sum( s[1][14] ),
					.cy( c[1][14] ));
assign sum[1] = s[1][14];

csa3 csa_s2_a0(
					.a( c[1][0] ),
					.b( c[1][1] ),
					.c( c[1][2] ),
					.sum( s[2][0] ),
					.cy( c[2][0] ));
csa3 csa_s2_a1(
					.a( s[2][0] ),
					.b( c[1][3] ),
					.c( c[1][4] ),
					.sum( s[2][1] ),
					.cy( c[2][1] ));
csa3 csa_s2_a2(
					.a( s[2][1] ),
					.b( c[1][5] ),
					.c( c[1][6] ),
					.sum( s[2][2] ),
					.cy( c[2][2] ));
csa3 csa_s2_a3(
					.a( s[2][2] ),
					.b( c[1][7] ),
					.c( c[1][8] ),
					.sum( s[2][3] ),
					.cy( c[2][3] ));
csa3 csa_s2_a4(
					.a( s[2][3] ),
					.b( c[1][9] ),
					.c( c[1][10] ),
					.sum( s[2][4] ),
					.cy( c[2][4] ));
csa3 csa_s2_a5(
					.a( s[2][4] ),
					.b( c[1][11] ),
					.c( c[1][12] ),
					.sum( s[2][5] ),
					.cy( c[2][5] ));
csa3 csa_s2_a6(
					.a( s[2][5] ),
					.b( c[1][13] ),
					.c( c[1][14] ),
					.sum( s[2][6] ),
					.cy( c[2][6] ));
assign sum[2] = s[2][6];

csa3 csa_s3_a0(
					.a( c[2][0] ),
					.b( c[2][1] ),
					.c( c[2][2] ),
					.sum( s[3][0] ),
					.cy( c[3][0] ));
csa3 csa_s3_a1(
					.a( s[3][0] ),
					.b( c[2][3] ),
					.c( c[2][4] ),
					.sum( s[3][1] ),
					.cy( c[3][1] ));
csa3 csa_s3_a2(
					.a( s[3][1] ),
					.b( c[2][5] ),
					.c( c[2][6] ),
					.sum( s[3][2] ),
					.cy( c[3][2] ));
assign sum[3] = s[3][2];

csa3 csa_s4_a0(
					.a( c[3][0] ),
					.b( c[3][1] ),
					.c( c[3][2] ),
					.sum( s[4][0] ),
					.cy( c[4][0] ));
assign sum[4] = s[4][0];

assign cy = c[4][0];


endmodule